
module top (

    //////////// CLOCK //////////
    input                       CLOCK_50,
    input                       CLOCK2_50,
    input                       CLOCK3_50,

    //////////// LED //////////
    output            [8:0]     LEDG,
    output           [17:0]     LEDR,

    //////////// KEY //////////
    input              [3:0]    KEY,

    //////////// SW //////////
    input             [17:0]    SW,

    //////////// SEG7 //////////
    output             [6:0]    HEX0,
    output             [6:0]    HEX1,
    output             [6:0]    HEX2,
    output             [6:0]    HEX3,
    output             [6:0]    HEX4,
    output             [6:0]    HEX5,
    output             [6:0]    HEX6,
    output             [6:0]    HEX7
);

//=======================================================
//  REG/WIRE declarations
//=======================================================

    /* 24 bit clock divider, converts 50MHz clock signal to 2.98Hz */
    logic [23:0] clkdiv;
    logic ledclk;
    assign ledclk = clkdiv[23];

    /* driver for LEDs */
    logic [25:0] leds;
    assign LEDR = leds[25:8];
    assign LEDG = leds[7:0];

    /* LED state register, 0 means going left, 1 means going right */
    logic ledstate;

    // --- define reset_n (active-low) and drive it from KEY[0] ---
    logic reset_n;
    assign reset_n = KEY[0];

//=======================================================
//  Behavioral coding
//=======================================================

    initial begin
        clkdiv = 26'h0;
        /* start at the far right, LEDG0 */
        leds = 26'b1;
        /* start out going to the left */
        ledstate = 1'b0;
    end

    always @(posedge CLOCK_50) begin
        /* drive the clock divider, every 2^26 cycles of CLOCK_50, the
        * top bit will roll over and give us a clock edge for clkdiv
        * */
        clkdiv <= clkdiv + 1;
    end

    always @(posedge ledclk) begin
        /* going left and we are at the far left, time to turn around */
        if ( (ledstate == 0) && (leds == 26'b10000000000000000000000000) ) begin
            ledstate <= 1;
            leds <= leds >> 1;

        /* going left and not at the far left, keep going */
        end else if (ledstate == 0) begin
            ledstate <= 0;
            leds <= leds << 1;

        /* going right and we are at the far right, turn around */
        end else if ( (ledstate == 1) && (leds == 26'b1) ) begin
            ledstate <= 0;
            leds <= leds << 1;

        /* going right, and we aren't at the far right */
        end else begin
            leds <= leds >> 1;
        end
    end
    
    logic        cpu_gpio_we;
    logic [31:0] cpu_gpio_wdata;
    logic [31:0] hex_data_reg;
    always_ff @(posedge CLOCK_50 or negedge KEY[0]) begin
        if (!KEY[0]) begin
            hex_data_reg <= 32'd0;
        end else if (cpu_gpio_we) begin
            hex_data_reg <= cpu_gpio_wdata;
        end
    end



    cpu u_cpu (
        .clk(CLOCK_50),                                                                                                                                                                                                  
        .rst_n      (reset_n),
        .io0_in     ({14'b0, SW}),   // zero-extend 18-bit switches
        .gpio_we    (cpu_gpio_we),   // strobe on csrrw HEX
        .gpio_wdata (cpu_gpio_wdata) // data written by csrrw HEX (rs1)
    );

    hexdriver disp0(.val(hex_data_reg[ 3: 0]), .HEX(HEX0)); // D0
    hexdriver disp1(.val(hex_data_reg[ 7: 4]), .HEX(HEX1)); // D1
    hexdriver disp2(.val(hex_data_reg[11: 8]), .HEX(HEX2)); // D2
    hexdriver disp3(.val(hex_data_reg[15:12]), .HEX(HEX3)); // D3
    hexdriver disp4(.val(hex_data_reg[19:16]), .HEX(HEX4)); // D4
    hexdriver disp5(.val(hex_data_reg[23:20]), .HEX(HEX5)); // D5
    hexdriver disp6(.val(hex_data_reg[27:24]), .HEX(HEX6)); // D6
    hexdriver disp7(.val(hex_data_reg[31:28]), .HEX(HEX7)); // D7

endmodule

