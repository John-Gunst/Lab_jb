
module top (

	//////////// CLOCK //////////
	input wire		          		CLOCK_50,
	input wire		          		CLOCK2_50,
	input wire		          		CLOCK3_50,

	//////////// KEY //////////
	input wire	     [3:0]		KEY,

	//////////// SW //////////
	input wire	    [17:0]		SW,

	//////////// SEG7 //////////
	output wire	     [6:0]		HEX0,
	output wire	     [6:0]		HEX1,
	output wire	     [6:0]		HEX2,
	output wire	     [6:0]		HEX3,
	output wire	     [6:0]		HEX4,
	output wire	     [6:0]		HEX5,
	output wire	     [6:0]		HEX6,
	output wire	     [6:0]		HEX7
);






//////////////////////////////////////////////////////////////////////////
// CPU board
//////////////////////////////////////////////////////////////////////////

	// internal wires for CPU to the board
	wire        cpu_rst;        // active high reset into cpu
	wire [31:0] cpu_gpio_in;    // CSR io0 (switches)
	wire [31:0] cpu_gpio_out;   // CSR io2 (hex display)
	wire        cpu_gpio_we;    // optional strobe when CPU writes io2

	// KEY[0] on DE2 is active-low. Convert to active-high reset for cpu.
	// if your cpu expects active low reset, pass KEY[0] directly instead.
	assign cpu_rst = ~KEY[0]; // press KEY0 -> cpu_rst = 1 (reset asserted)

	// zero extend SW into 32-bit CSR input
	assign cpu_gpio_in = {14'd0, SW}; // adjust if your SW width differs

	// instantiate the CPU
	cpu u_cpu (
	    .clk      (CLOCK_50),    // board clock
	    .rst      (cpu_rst),     // cpu reset
	    .gpio_in  (cpu_gpio_in),
	    .gpio_out (cpu_gpio_out)
	    //.gpio_we  (cpu_gpio_we)
	);

	// instantiate hexdrivers: map packed 32-bit cpu_gpio_out -> HEX0..HEX7
	// LSB 4bits -> HEX0, next 4bits -> HEX1, etc.
	hexdriver hd0 (.val(cpu_gpio_out[3:0]),   .HEX(HEX0));
	hexdriver hd1 (.val(cpu_gpio_out[7:4]),   .HEX(HEX1));
	hexdriver hd2 (.val(cpu_gpio_out[11:8]),  .HEX(HEX2));
	hexdriver hd3 (.val(cpu_gpio_out[15:12]), .HEX(HEX3));
	hexdriver hd4 (.val(cpu_gpio_out[19:16]), .HEX(HEX4));
	hexdriver hd5 (.val(cpu_gpio_out[23:20]), .HEX(HEX5));
	hexdriver hd6 (.val(cpu_gpio_out[27:24]), .HEX(HEX6));
	hexdriver hd7 (.val(cpu_gpio_out[31:28]), .HEX(HEX7));

	// optional debug: light an LED when cpu writes to the HEX CSR
	// assign LEDR[0] = cpu_gpio_we;
endmodule
